/*************************************************

 Copyright: NUDT_CoreLight

 File name: upsp_pkg.sv

 Author: NUDT_CoreLight

 Date: 2021-04-13


 Description:


 **************************************************/

package upsp_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "upsp_trans.svh"

`include "upsp_driver.svh"
`include "upsp_monitor.svh"
`include "upsp_sqr.svh"

`include "upsp_ostream_modifier.svh"

`include "upsp_agent.svh"

endpackage