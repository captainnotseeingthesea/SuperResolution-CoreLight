/*************************************************

 Copyright: NUDT_CoreLight

 File name: ifs.sv

 Author: NUDT_CoreLight

 Date: 2021-04-15


 Description:

 SV interfaces for verification.

 **************************************************/


`include "axi_lite_if.svh"

`include "axi_stream_if.svh"

`include "upsp_if.svh"

`include "ac_if.svh"

