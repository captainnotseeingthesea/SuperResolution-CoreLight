/*************************************************

 Copyright: NUDT_CoreLight

 File name: axi_lite_pkg.sv

 Author: NUDT_CoreLight

 Date: 2021-04-13


 Description:


 **************************************************/

package axi_lite_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "axi_lite_trans.svh"

`include "m_axi_lite_driver.svh"
`include "m_axi_lite_sqr.svh"
`include "m_axi_lite_agent.svh"

endpackage