/*************************************************

 Copyright: NUDT_CoreLight

 File name: duts.sv

 Author: NUDT_CoreLight

 Date: 2021-04-06


 Description:

 DUTs

 **************************************************/

`include "ac_crf_top.svh"

`include "bcci_ip_top.svh"