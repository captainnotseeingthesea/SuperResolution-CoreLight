/*************************************************

 Copyright: NUDT_CoreLight

 File name: utils_pkg.sv

 Author: NUDT_CoreLight

 Date: 2021-04-14


 Description:

 Usefult utilities 

 **************************************************/

package utils_pkg;

    string utils_path = "";

`include "bmp.svh"


endpackage